module ISERDESE2 #(
   parameter         DATA_RATE           = "DDR",
   parameter integer DATA_WIDTH          = 4,
   parameter         DYN_CLKDIV_INV_EN   = "FALSE",
   parameter         DYN_CLK_INV_EN      = "FALSE",
   parameter [0:0]   INIT_Q1             = 1'b0,
   parameter [0:0]   INIT_Q2             = 1'b0,
   parameter [0:0]   INIT_Q3             = 1'b0,
   parameter [0:0]   INIT_Q4             = 1'b0,
   parameter         INTERFACE_TYPE      = "MEMORY",
   parameter         IOBDELAY            = "NONE",
   parameter [0:0]   IS_CLKB_INVERTED    = 1'b0,
   parameter [0:0]   IS_CLKDIVP_INVERTED = 1'b0,
   parameter [0:0]   IS_CLKDIV_INVERTED  = 1'b0,
   parameter [0:0]   IS_CLK_INVERTED     = 1'b0,
   parameter [0:0]   IS_D_INVERTED       = 1'b0,
   parameter [0:0]   IS_OCLKB_INVERTED   = 1'b0,
   parameter [0:0]   IS_OCLK_INVERTED    = 1'b0,
   parameter integer NUM_CE              = 2,
   parameter         OFB_USED            = "FALSE",
   parameter         SERDES_MODE         = "MASTER",
   parameter [0:0]   SRVAL_Q1            = 1'b0,
   parameter [0:0]   SRVAL_Q2            = 1'b0,
   parameter [0:0]   SRVAL_Q3            = 1'b0,
   parameter [0:0]   SRVAL_Q4            = 1'b0
)(
   output O,
   output Q1,
   output Q2,
   output Q3,
   output Q4,
   output Q5,
   output Q6,
   output Q7,
   output Q8,
   output SHIFTOUT1,
   output SHIFTOUT2,

   input  BITSLIP,
   input  CE1,
   input  CE2,
   input  CLK,
   input  CLKB,
   input  CLKDIV,
   input  CLKDIVP,
   input  D,
   input  DDLY,
   input  DYNCLKDIVSEL,
   input  DYNCLKSEL,
   input  OCLK,
   input  OCLKB,
   input  OFB,
   input  RST,
   input  SHIFTIN1,
   input  SHIFTIN2
);
endmodule: ISERDESE2
