//======================================================================== 
// openeye-CamSI * NLnet-sponsored open-source core for Camera I/F with ISP
//------------------------------------------------------------------------
//                   Copyright (C) 2024 Chili.CHIPS*ba
// 
// Redistribution and use in source and binary forms, with or without 
// modification, are permitted provided that the following conditions 
// are met:
//
// 1. Redistributions of source code must retain the above copyright 
// notice, this list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright 
// notice, this list of conditions and the following disclaimer in the 
// documentation and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its 
// contributors may be used to endorse or promote products derived
// from this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS 
// IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED 
// TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A 
// PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT 
// HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, 
// SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT 
// LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, 
// DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY 
// THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT 
// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE 
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
//              https://opensource.org/license/bsd-3-clause
//------------------------------------------------------------------------
// Designers  : Armin Zunic, Isam Vrce
// Description: AXI Streaming (Data Plane) interface. For more, see:
//               https://zipcpu.com/doc/axi-stream.pdf
//========================================================================

interface axis_if #(
   parameter DWIDTH = 64,         // allowed values are 64, 128, 256, 512, 1024 
   parameter KWIDTH = DWIDTH / 8, // width of KEEP bus: DMA=DWIDTH/8
   parameter UWIDTH = 1           // width of TUSER bus
); 

   logic              TREADY;
   logic              TVALID;
   logic [DWIDTH-1:0] TDATA;
   logic [KWIDTH-1:0] TKEEP;
   logic              TLAST;

   logic [UWIDTH-1:0] TUSER;
   

  //---------------------------------------- 
  // MASTER side
  //---------------------------------------- 
   modport MASTER (
      input  TREADY,

      output TVALID,
      output TDATA,
      output TKEEP,
      output TLAST,

      output TUSER
   );


  //---------------------------------------- 
  // SLAVE side
  //---------------------------------------- 
   modport SLAVE (
      output TREADY,

      input  TVALID,
      input  TDATA,
      input  TKEEP,
      input  TLAST,

      input  TUSER
   );

endinterface: axis_if

/*
-----------------------------------------------------------------------------
Version History:
-----------------------------------------------------------------------------
 2024/01/15 AZ: initial creation    

*/
